grammar edu:umn:cs:melt:exts:ableC:checkTaggedUnion;

exports edu:umn:cs:melt:exts:ableC:checkTaggedUnion:abstractsyntax;

