grammar determinism;

import edu:umn:cs:melt:ableC:host;

copper_mda testStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:check;
  edu:umn:cs:melt:exts:ableC:checkTaggedUnion;
}

