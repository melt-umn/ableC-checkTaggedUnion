grammar edu:umn:cs:melt:exts:ableC:taggedUnion;

exports edu:umn:cs:melt:exts:ableC:taggedUnion:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:taggedUnion:concretesyntax;

